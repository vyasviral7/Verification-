module viral()

$display ("VIRAL VIRAL");

endmodule
